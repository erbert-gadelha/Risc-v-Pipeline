`timescale 1ns / 1ps

module Controller (
    //Input
    input logic [6:0] Opcode,
    //7-bit opcode field from the instruction

    //Outputs
    output logic ALUSrc,
    //0: The second ALU operand comes from the second register file output (Read data 2); 
    //1: The second ALU operand is the sign-extended, lower 16 bits of the instruction.
    output logic MemtoReg,
    //0: The value fed to the register Write data input comes from the ALU.
    //1: The value fed to the register Write data input comes from the data memory.
    output logic RegWrite, //The register on the Write register input is written with the value on the Write data input 
    output logic MemRead,  //Data memory contents designated by the address input are put on the Read data output
    output logic MemWrite, //Data memory contents designated by the address input are replaced by the value on the Write data input.
    output logic [1:0] ALUOp,  //00: LW/SW; 01:Branch; 10: Rtype
    output logic Branch  //0: branch is not taken; 1: branch is taken
);

  logic [6:0] R_TYPE, LW, SW, BR;

  assign R_TYPE    = 7'b0110011;  // [R_TYPE] add,and (diferenciar pelo campo funct3 e funct7)
  assign LOAD      = 7'b0000011;  // [I-TYPE] LB, LH, LW, LBU, LHU
  assign STORE     = 7'b0100011;  // [S-TYPE] SB, SH, SW
  assign BRANCH    = 7'b1100011;  // [B-TYPE] BEQ, BNE, BLT, BGE, ...
  assign IMMEDIATE = 7'b0010011;  // [I-TYPE] ADDI, XORI, ... 
  assign JAL       = 7'b1101111;  // [J-TYPE]
  assign JALR      = 7'b1101111;  // [J-TYPE]
  assign LUI       = 7'b1101111;  // [U-TYPE]
  assign SYSCALL   = 7'b1110011;  // HALT

  assign ALUSrc   = (Opcode == LOAD || Opcode == STORE);
  assign MemtoReg = (Opcode == LOAD);
  assign RegWrite = (Opcode == R_TYPE || Opcode == LOAD);
  assign MemRead  = (Opcode == LOAD);
  assign MemWrite = (Opcode == STORE);
  assign ALUOp[0] = (Opcode == BRANCH);
  assign ALUOp[1] = (Opcode == R_TYPE);
  assign Branch   = (Opcode == BRANCH);

endmodule
